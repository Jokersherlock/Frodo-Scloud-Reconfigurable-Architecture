`timescale 1ns / 1ns

// `define USE_IP

// `define PRINT_RAM